module NB_DIGITAL_TOP_tb();
  /*autowire*/
  /*autoreginput*/


  NB_DIGITAL_TOP nb_digital_top
  (/*autoinst*/);  

endmodule
